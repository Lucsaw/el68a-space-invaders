library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

library work;
use work.spaceInvadersConstants.all;

entity spaceInvaders is
	port (
		clk, rst                          : in std_logic
	);
end spaceInvaders;

architecture aSpaceInvaders of spaceInvaders is
  

begin

  
  
end architecture aSpaceInvaders;