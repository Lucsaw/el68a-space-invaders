library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity spaceInvaders is
  port (
    clock   : in std_logic;
    rst     : in std_logic
  );
end spaceInvaders;

architecture aSpaceInvaders of spaceInvaders is
  
begin
  
  
  
end architecture aSpaceInvaders;